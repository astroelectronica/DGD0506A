.title KiCad schematic
.include "C:/AE/DGD0506A/DGD0506A.spice.txt"
.include "C:/AE/DGD0506A/DMN6017SK3.spice.txt"
.include "C:/AE/DGD0506A/c2012x7r2a104k125ae_p.mod"
.include "C:/AE/DGD0506A/c3216x6s2a106k160ac_p.mod"
.include "C:/AE/DGD0506A/cga4j3x7s2a105k125ae_p.mod"
XU2 VCC 0 C2012X7R2A104K125AE_p
R1 0 /DT {RDT}
R4 /ENABLE VCC {RPU}
XU1 VCC /VB /HO /OUTPUT unconnected-_U1-NC-Pad5_ /DT /ENABLE /INPUT 0 /LO dgd0506a
V3 /INPUT 0 DC PULSE(0 {VPUL} {DELAY} {TR} {TF} {DUTY} {CYCLE}) 
R5 0 /OUTPUT {RLOAD}
XQ1 VBUS /GHO /OUTPUT DMN6017SK3
XQ2 /OUTPUT /GLO 0 DMN6017SK3
R3 /GHO /HO {RHO}
R2 /GLO /LO {RLO}
XU3 /VB /OUTPUT CGA4J3X7S2A105K125AE_p
XU4 VBUS 0 C3216X6S2A106K160AC_p
V1 VCC 0 DC {VCC} 
V2 VBUS 0 DC {VBUS} 
.end
