.title KiCad schematic
.include "C:/AE/DGD0506A/DGD0506A.spice.txt"
.include "C:/AE/DGD0506A/DMN6017SK3.spice.txt"
R1 0 /DT {RDT}
XU1 VCC /VB /HO /OUTPUT unconnected-_U1-NC-Pad5_ /DT /ENABLE /INPUT 0 /LO dgd0506a
R4 /ENABLE VCC {RPU}
C1 VCC 0 100n
V3 /INPUT 0 DC PULSE(0 {VPUL} {DELAY} {TR} {TF} {DUTY} {CYCLE}) 
C3 VBUS 0 10u
C2 /VB /OUTPUT 100n
R3 /GHO /HO {RHO}
R2 /GLO /LO {RLO}
XQ2 /OUTPUT /GLO 0 DMN6017SK3
XQ1 VBUS /GHO /OUTPUT DMN6017SK3
R5 0 /OUTPUT {RLOAD}
V2 VBUS 0 DC {VBUS} 
V1 VCC 0 DC {VCC} 
.end
